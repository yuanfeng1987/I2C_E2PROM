// State definition
`define Idle 3'b000
`define Start 3'b001
`define Chip_Addr_Send 3'b010
`define Reg_Addr_Send 3'b011
`define Data_Send 3'b100
`define Data_Rcv 3'b101
`define Stop 3'b110

// flag definition 
// whether I2C module is enabled or not: 
`define I2C_disabled 1'b0
`define I2C_Enabled 1'b1
//I2C module read or write enabled :i_R_W
`define Read_Enabled 1'b1
`define Wrt_Enabled 1'b0
// The receiving or sending data is finished or not : 
`define Data_RS_Done 1'b0
`define Data_RS_NotDone 1'b1
// The E2PROM current addr is the required addr
`define Read_Setting_Done 1'b1
`define Read_Setting_NotDone 1'b0
// The clock time reached the preset value, the current action is done
`define Time_Expired  1'b0
`define Time_NotExpired  1'b1
// whether fault occurs during current state:
`define Err_Yes 1'b1
`define Err_No  1'b0

// timer expiraion value definition
`define Start_Timer 8'b0010_1000
`define Start_Timer_Ph1 8'b0000_1111
`define Start_Timer_Ph2 8'b0001_1001

`define RS_Data_Timer 8'b1110_0001

`define Stop_Timer 8'b0010_1000
`define Stop_Timer_Ph1 8'b0000_1111
`define Stop_Timer_Ph2 8'b0001_1001

module State_Transfer(input wire i_RST_n,				  // system reset
							 input wire i_clk10MHz,			  // clock generated by system PLL
							 input wire i_I2C_Enable_Flag,			  // I2C enbbled by CPU
							 input wire i_R_W,				  // Read or write icon: 1, read; 0, write
							 input wire i_Num_Remain,		  // the number of sending or received data: 0, finished; 1, not finished
							 input wire i_Read_Setting_Flag,     // the E2PROM read is enabled or not: 1, enabled; 0, not enabled.
							 input wire i_Timer_Flag,            // current state time during expired or not: 0, expired; 1, not expired 
							 input wire i_Err_Flag,              // sending or receiving error occurs
							 
							 output reg [2:0] Current_State);
	reg [2:0] Next_state;
	
	
	always @(posedge i_clk10MHz or negedge i_RST_n)    // transfer to next state
	begin 
		if(!i_RST_n)
			begin
				Current_State<=`Idle;
			end
		else
			begin
				Current_State<=Next_state;
			end
	end
	
	always @(*)
	begin
		if(!i_RST_n)
		begin
			Next_state<=`Idle;
		end
		else 
			case (Current_State)
			`Idle: begin
					if(i_I2C_Enable_Flag==`I2C_Enabled)
						Next_state<=`Start;
					else
						Next_state<=`Idle;
					end
			`Start: begin
					if (i_Timer_Flag==`Time_NotExpired)
						Next_state<=`Start;
					else
						Next_state<=`Chip_Addr_Send;
					end
			`Chip_Addr_Send: begin
					if (i_Timer_Flag==`Time_NotExpired) // not expired
						Next_state<=`Chip_Addr_Send;
					else if ((i_R_W==`Read_Enabled)&(i_Read_Setting_Flag==`Read_Setting_Done))
						Next_state<=`Data_Rcv;
					else
						Next_state<=`Reg_Addr_Send ;
					end
			`Data_Rcv: begin
					if (i_Timer_Flag==`Time_NotExpired)
						Next_state<=`Data_Rcv;
					else if (i_Num_Remain==`Data_RS_NotDone)
						Next_state<=`Data_Rcv;	
					else
						Next_state<=`Stop;
			      end
			`Reg_Addr_Send: begin
					if (i_Timer_Flag==`Time_NotExpired)
						Next_state<=`Reg_Addr_Send;
					else if (i_R_W==`Read_Enabled)      // whether setting flag should be enabled ?
						Next_state<=`Start;
					else
					   Next_state<=`Data_Send;
					end
			`Data_Send: begin
					if (i_Timer_Flag==`Time_NotExpired)
						Next_state<=`Data_Send;
					else if(i_Num_Remain==`Data_RS_NotDone)
						Next_state<=`Data_Send;
					else
						Next_state<=`Stop;
					end
			`Stop: begin
					if (i_Timer_Flag==`Time_NotExpired)
						Next_state<=`Stop;
					else
						Next_state<=`Idle;
					end
			default:
						Next_state<=`Idle;
			endcase
	end
	
endmodule